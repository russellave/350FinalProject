module modulo(score,out);
input [9:0] score;
output [20:0] out;

wire [5:0] hundred;
wire [5:0] ten;
wire [5:0] one;
assign hundred = score % 100;
assign ten = score % 10;
assign one = score % 1;
assign out [6:0] = 	({7{(one == 5'h0)}} & 7'b1000000) |
		({7{(one == 6'h1)}} & 7'b1111001) |
		({7{(one == 6'h2)}} & 7'b0100100) |
		({7{(one == 6'h3)}} & 7'b0110000) |
		({7{(one == 6'h4)}} & 7'b0011001) |
		({7{(one == 6'h5)}} & 7'b0010010) |
		({7{(one == 6'h6)}} & 7'b0000010) |
		({7{(one == 6'h7)}} & 7'b1111000) |
		({7{(one == 6'h8)}} & 7'b0000000) |
		({7{(one == 6'h9)}} & 7'b0010000);
assign out [13:7] = 	({7{(ten == 5'h0)}} & 7'b1000000) |
		({7{(ten == 6'h1)}} & 7'b1111001) |
		({7{(ten == 6'h2)}} & 7'b0100100) |
		({7{(ten == 6'h3)}} & 7'b0110000) |
		({7{(ten == 6'h4)}} & 7'b0011001) |
		({7{(ten == 6'h5)}} & 7'b0010010) |
		({7{(ten == 6'h6)}} & 7'b0000010) |
		({7{(ten == 6'h7)}} & 7'b1111000) |
		({7{(ten == 6'h8)}} & 7'b0000000) |
		({7{(ten == 6'h9)}} & 7'b0010000);
assign out [20:14] = 	({7{(hundred == 5'h0)}} & 7'b1000000) |
		({7{(hundred == 6'h1)}} & 7'b1111001) |
		({7{(hundred == 6'h2)}} & 7'b0100100) |
		({7{(hundred == 6'h3)}} & 7'b0110000) |
		({7{(hundred == 6'h4)}} & 7'b0011001) |
		({7{(hundred == 6'h5)}} & 7'b0010010) |
		({7{(hundred == 6'h6)}} & 7'b0000010) |
		({7{(hundred == 6'h7)}} & 7'b1111000) |
		({7{(hundred == 6'h8)}} & 7'b0000000) |
		({7{(hundred == 6'h9)}} & 7'b0010000);	
endmodule