module skeleton(resetn, 
	ps2_clock, ps2_data, 										// ps2 related I/O
	debug_data_in, debug_addr, leds, 						// extra debugging ports
	lcd_data, lcd_rw, lcd_en, lcd_rs, lcd_on, lcd_blon,// LCD info
	seg1, seg2, seg3, seg4, seg5, seg6, seg7, seg8,		// seven segements
	VGA_CLK,   														//	VGA Clock
	VGA_HS,															//	VGA H_SYNC
	VGA_VS,															//	VGA V_SYNC
	VGA_BLANK,														//	VGA BLANK
	VGA_SYNC,														//	VGA SYNC
	VGA_R,   														//	VGA Red[9:0]
	VGA_G,	 														//	VGA Green[9:0]
	VGA_B,															//	VGA Blue[9:0]
	CLOCK_50, sensor_input, out_final, final_sensor_output, controller, controller_output, save_signal, load_signal, sensor_input_out, state_load_out, counter, CLOCK_27,
	KEY, SW, AUD_ADCDAT, AUD_BCLK, AUD_ADCLRCK, AUD_DACLRCK, I2C_SDAT, AUD_XCK, AUD_DACDAT, I2C_SCLK, scoreconverted);  													// 50 MHz clock
		
	////////////////////////	VGA	////////////////////////////
	output			VGA_CLK;   				//	VGA Clock
	output			VGA_HS;					//	VGA H_SYNC
	output			VGA_VS;					//	VGA V_SYNC
	output			VGA_BLANK;				//	VGA BLANK
	output			VGA_SYNC;				//	VGA SYNC
	output	[7:0]	VGA_R;   				//	VGA Red[9:0]
	output	[7:0]	VGA_G;	 				//	VGA Green[9:0]
	output	[7:0]	VGA_B;   				//	VGA Blue[9:0]
	input				CLOCK_50;

	////////////////////////	PS2	////////////////////////////
	input 			resetn;
	inout 			ps2_data, ps2_clock;
	
	////////////////////////	LCD and Seven Segment	////////////////////////////
	output 			   lcd_rw, lcd_en, lcd_rs, lcd_on, lcd_blon;
	output 	[7:0] 	leds, lcd_data;
	output 	[6:0] 	seg1, seg2, seg3, seg4, seg5, seg6, seg7, seg8;
	output 	[31:0] 	debug_data_in;
	output   [11:0]   debug_addr;
	output [20:0] scoreconverted;
	
	
	
	
	wire			 clock;
	wire			 lcd_write_en;
	wire 	[31:0] lcd_write_data;
	wire	[7:0]	 ps2_key_data;
	wire			 ps2_key_pressed;
	wire	[7:0]	 ps2_out;	
	
	//Final Project 
	
	input [31:0] sensor_input; //only first (lsb) 24 bits matter. goes to vga controller and processor (address 0)
	output [31:0] sensor_input_out; 
	assign sensor_input_out = sensor_input; 
	//output processor
	output [31:0] final_sensor_output; //only first 3 bits matter. which light to turn on (address 1)
	
	input [31:0] controller; //only first 3 bits matter. goes to processor (address 2)
	output [31:0] controller_output; 
	
	assign controller_output = controller; 

	//output vga
	wire [31:0] sensor_input_to_save; 
	output [31:0] save_signal; 
	output [31:0] load_signal; 
	output [2:0] state_load_out; 
	output [31:0] counter; 
	wire [31:0] sensor_output; 
	wire [31:0] adjusted_sensor_output; 
	wire [31:0] screen_out; 
	wire [31:0] out_game; 
	// clock divider (by 5, i.e., 10 MHz)
	pll div(CLOCK_50,inclock);
	assign clock = CLOCK_50;
	
	// UNCOMMENT FOLLOWING LINE AND COMMENT ABOVE LINE TO RUN AT 50 MHz
//   assign clock = inclock;
	
	// your processor
//	processor_skeleton myprocessor(clock, ~resetn, sensor_input, sensor_output, save_signal, load_signal, counter/*ps2_key_pressed, ps2_out, lcd_write_en, lcd_write_data,*/);
	wire [31:0] not_controller; 
	not not1(not_controller[0], controller[0]);
	not not2(not_controller[1], controller[1]);
	not not3(not_controller[2], controller[2]);
	not not4(not_controller[3], controller[3]);
	processor_skeleton_alt myprocessor_alt(clock, ~resetn, sensor_input, sensor_output, not_controller, screen_out/*ps2_key_pressed, ps2_out, lcd_write_en, lcd_write_data,*/ );
	
	// keyboard controller
	PS2_Interface myps2(clock, resetn, ps2_clock, ps2_data, ps2_key_data, ps2_key_pressed, ps2_out);
	
	// lcd controller
	lcd mylcd(clock, ~resetn, 1'b1, ps2_out, lcd_data, lcd_rw, lcd_en, lcd_rs, lcd_on, lcd_blon);
	
	// example for sending ps2 data to the first two seven segment displays
	Hexadecimal_To_Seven_Segment hex1(ps2_out[3:0], seg1);
	Hexadecimal_To_Seven_Segment hex2(ps2_out[7:4], seg2);
	
	// the other seven segment displays are currently set to 0
	Hexadecimal_To_Seven_Segment hex3(4'b0, seg3);
	Hexadecimal_To_Seven_Segment hex4(4'b0, seg4);
	Hexadecimal_To_Seven_Segment hex5(4'b0, seg5);
	Hexadecimal_To_Seven_Segment hex6(4'b0, seg6);
	Hexadecimal_To_Seven_Segment hex7(4'b0, seg7);
	Hexadecimal_To_Seven_Segment hex8(4'b0, seg8);
	
	// some LEDs that you could use for debugging if you wanted
	assign leds = 8'b00101011;
	
//   or or_pad1(adjusted_sensor_output[0], ~sensor_output[0], ~sensor_output[1], ~sensor_output[2], ~sensor_output[3], ~sensor_output[4]);
//	or or_pad2(adjusted_sensor_output[1], ~sensor_output[5], ~sensor_output[6], ~sensor_output[7], ~sensor_output[8], ~sensor_output[9]);
//	or or_pad3(adjusted_sensor_output[2], ~sensor_output[14], ~sensor_output[13], ~sensor_output[12], ~sensor_output[11], ~sensor_output[10]);
//	
		
	// VGA
	Reset_Delay			r0	(.iCLK(CLOCK_50),.oRESET(DLY_RST)	);
	VGA_Audio_PLL 		p1	(.areset(~DLY_RST),.inclk0(CLOCK_50),.c0(VGA_CTRL_CLK),.c1(AUD_CTRL_CLK),.c2(VGA_CLK)	);
//	vga_controller vga_ins(.iRST_n(DLY_RST),
//								 .iVGA_CLK(VGA_CLK),
//								 .oBLANK_n(VGA_BLANK),
//								 .oHS(VGA_HS),
//								 .oVS(VGA_VS),
//								 .b_data(VGA_B),
//								 .g_data(VGA_G),
//								 .r_data(VGA_R), 
//								 .sensor_input(sensor_input), //input
//								 .sensor_output_adjusted(adjusted_sensor_output), //input
//								 .controller(controller), //input
//								 .sensor_input_to_save(sensor_input_to_save), //output to processor
//								 .save_signal(save_signal), //output to processor
//								 .load_signal(load_signal), 
//								 .state_load_out(state_load_out), 
//								 .load_counter(counter), //output to processor
//								 .final_out_dummy(final_sensor_output)); 

	vga_controller_alt vga_ins_alt(.iRST_n(DLY_RST),
								 .iVGA_CLK(VGA_CLK),
								 .oBLANK_n(VGA_BLANK),
								 .oHS(VGA_HS),
								 .oVS(VGA_VS),
								 .b_data(VGA_B),
								 .g_data(VGA_G),
								 .r_data(VGA_R), 
							 .sensor_input(sensor_input), 
							 .screen(screen_out),
							 .out_game(out_game),
							 .scoreconverted(scoreconverted));
	wire case_game; 
	output [31:0] out_final; 
	assign out_final = out_game; 
//	or or_out_game_not_zero(out_game[0], out_game[1], out_game[2], out_game[3], out_game[4], out_game[5]); 
//	assign out_final = case_game ? out_game : sensor_output;  
	
	
	wire game_over; 
	assign game_over = 1'b0; 
	
	input				CLOCK_27;  
	input		[3:0]	KEY;
	input		[3:0]	SW;

	input				AUD_ADCDAT;

	// Bidirectionals
	inout				AUD_BCLK;
	inout				AUD_ADCLRCK;
	inout				AUD_DACLRCK;

	inout				I2C_SDAT;

	// Outputs
	output				AUD_XCK;
	output				AUD_DACDAT;

	output				I2C_SCLK;
	DE2_Audio_Example audio_inst (
	.game_over(game_over),
	// Inputs
	.CLOCK_50(CLOCK_50),
	.AUD_ADCDAT(AUD_ADCDAT),
	.KEY(KEY),
	
	// Bidirectionals
	.AUD_BCLK(AUD_BCLK),
	.AUD_ADCLRCK(AUD_ADCLRCK),
	.AUD_DACLRCK(AUD_DACLRCK),

	.I2C_SDAT(I2C_SDAT),

	// Outputs
	.AUD_XCK(AUD_XCK),
	.AUD_DACDAT(AUD_DACDAT),

	.I2C_SCLK(I2C_SCLK)
	);
	
endmodule
